module controller(

);

// forwarding

// jump

// memeory hazard

endmodule